`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2017/12/12 11:26:03
// Design Name: 
// Module Name: hilo_reg
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module hilo_reg(
	input  wire clk,rst,we,
	input wire diven,
	input wire [5:0] alucontrol,
	input wire [63:0] div_result,
	input  wire [31:0] hi_i,lo_i,
	output wire [31:0] hi_o,lo_o
    );
	
	reg [31:0] hi, lo;
	always @(posedge clk) begin
		if(rst) begin
			hi <= 0;
			lo <= 0;
		end else if (we) begin
		    if(diven)begin
		        hi<=div_result[63:32];
		        lo<=div_result[31:0];
		    end else if (alucontrol==`MTHI_CONTROL | alucontrol==`MTLO_CONTROL
		     | alucontrol==`MULT_CONTROL | alucontrol==`MULTU_CONTROL) begin
			     hi <= hi_i;
			     lo <= lo_i;
			end
		end
	end

	assign hi_o = hi;
	assign lo_o = lo;
endmodule

`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2024/01/09 17:31:41
// Design Name: 
// Module Name: mips_top
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module mips_core(
    input wire clk,
    input wire resetn,  //low active
    input wire [5:0] ext_int,

    //instr
    output wire inst_req,
    output wire inst_wr,
    output wire [1:0] inst_size,
    output wire [31:0] inst_addr,
    output wire [31:0] inst_wdata,
    input wire inst_addr_ok,
    input wire inst_data_ok,
    input wire [31:0] inst_rdata,

    //data
    output wire data_req,
    output wire data_wr,
    output wire [1:0] data_size,
    output wire [31:0] data_addr,
    output wire [31:0] data_wdata,
    input wire data_addr_ok,
    input wire data_data_ok,
    input wire [31:0] data_rdata,

    //debug
    output wire [31:0] debug_wb_pc,
    output wire [3:0] debug_wb_rf_wen ,
    output wire [4:0] debug_wb_rf_wnum ,
    output wire [31:0] debug_wb_rf_wdata
);

	wire [31:0] instr;
	wire [3:0] memwrite;
	wire [31:0] aluoutM, writedata, readdataM,result,pcW;
	wire regwrite;
	wire [4:0] writereg;
	
	//sram
    wire i_stall,d_stall,longest_stall;
    wire [31:0] inst_sram_rdata;
    wire [31:0] inst_sram_addr ;
    wire inst_sram_en,data_sram_en;
	    
    mips mips(
        .clk(clk),
        .rst(resetn),
        .ext_int(ext_int),
        //instr
        // .inst_en(inst_en),
        .pcF(inst_sram_addr),                    //pcF
        .instrF(inst_sram_rdata),              //instrF
        //data
        // .data_en(data_en),
        .aluoutM(aluoutM),
        .writedataM(writedata),
        .readdataM(readdataM),
        .memwriteM(memwrite),
        .pcW(pcW),
        .resultW(result),
        .writeregW(writereg),
        .regwriteW(regwrite),
        .data_sram_en(data_sram_en),
        .inst_enF(inst_sram_en),
        .i_stall(i_stall),.d_stall(d_stall),
        .longest_stall(longest_stall)
    );

    assign debug_wb_pc = pcW;
    assign debug_wb_rf_wen ={4{regwrite}};
    assign debug_wb_rf_wnum = writereg;
    assign debug_wb_rf_wdata = result;

        //inst sram to sram-like
    i_sram_like i_sram_to_sram_like(
        .clk(clk), .rst(resetn),
        //sram
        .inst_sram_en(inst_sram_en),
        .inst_sram_addr(inst_sram_addr),
        .inst_sram_rdata(inst_sram_rdata),
        .i_stall(i_stall),
        .longest_stall(longest_stall),
        //sram like
        .inst_req(inst_req), 
        .inst_wr(inst_wr),
        .inst_size(inst_size),
        .inst_addr(inst_addr),   
        .inst_wdata(inst_wdata),
        .inst_addr_ok(inst_addr_ok),
        .inst_data_ok(inst_data_ok),
        .inst_rdata(inst_rdata)    
    );

    //data sram to sram-like
    d_sram_like d_sram_to_sram_like(
        .clk(clk), .rst(resetn),
        //sram
        .data_sram_en(data_sram_en),
        .data_sram_addr(aluoutM),
        .data_sram_rdata(readdataM),
        .data_sram_wen(memwrite),
        .data_sram_wdata(writedata),
        .d_stall(d_stall),
        .longest_stall(longest_stall),
        //sram like
        .data_req(data_req),    
        .data_wr(data_wr),
        .data_size(data_size),
        .data_addr(data_addr),   
        .data_wdata(data_wdata),
        .data_addr_ok(data_addr_ok),
        .data_data_ok(data_data_ok),
        .data_rdata(data_rdata)
    );
    
    //ascii
    instdec instdec(
        .instr(inst_sram_rdata)
    );

endmodule
